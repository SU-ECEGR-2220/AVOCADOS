--------------------------------------------------------------------------------
--
-- LAB #4
--
--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity fulladder is
    port (a : in std_logic;
          b : in std_logic;
          cin : in std_logic;
          sum : out std_logic;
          carry : out std_logic
         );
end fulladder;

architecture addlike of fulladder is
begin
  sum   <= a xor b xor cin; 
  carry <= (a and b) or (a and cin) or (b and cin); 
end architecture addlike;

--------------------------------------------------------------------------------

Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity adder_subtracter is
	port(	datain_a: in std_logic_vector(31 downto 0);
		datain_b: in std_logic_vector(31 downto 0);
		add_sub: in std_logic;
		dataout: out std_logic_vector(31 downto 0);
		co: out std_logic);
end entity adder_subtracter;

architecture calc of adder_subtracter is
	-- insert component
	component fulladder
		port (a: in std_logic;
		      b: in std_logic;
		      cin: in std_logic;
		      sum: out std_logic;
		      carry: out std_logic);
	end component;

	-- creating signal for data of b and carries
	signal db: std_logic_vector(31 downto 0);
	signal c: std_logic_vector(32 downto 0);

begin
	with add_sub select
		db <= 	datain_b when '0',  		-- db = B when add
			not(datain_b) when others;	-- db = -B when subtract
	c(0) <= add_sub;
	co <= c(32); -- data in 32th-bit-carry is carryout
 
	-- create loop to run fulladder component
	add32: for i in 0 to 31 generate
	f: fulladder port map (datain_a(i),db(i),c(i),dataout(i),c(i+1));
	end generate;

	
end architecture calc;


--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity shift_register is
	port(	datain: in std_logic_vector(31 downto 0);
	   	dir: in std_logic;
		shamt:	in std_logic_vector(4 downto 0);
		dataout: out std_logic_vector(31 downto 0));
end entity shift_register;

architecture shifter of shift_register is
	
begin
	-- insert code here.
	with dir & shamt select
		dataout <= datain(30 downto 0) & '0'   when "000001",
			   datain(29 downto 0) & "00"  when "000010",
			   datain(28 downto 0) & "000" when "000011",

			   '0'   & datain(31 downto 1) when "100001",
			   "00"  & datain(31 downto 2) when "100010",
			   "000" & datain(31 downto 3) when "100011",
			   datain(31 downto 0) when others;

end architecture shifter;


--------------------------------------------------------------------------------

Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity ALU is
	Port(	DataIn1: in std_logic_vector(31 downto 0);
		DataIn2: in std_logic_vector(31 downto 0);
		ALUCtrl: in std_logic_vector(4 downto 0);
		Zero: out std_logic;
		ALUResult: out std_logic_vector(31 downto 0) );
end entity ALU;

architecture ALU_Arch of ALU is
	signal addsub_result: std_logic_vector(31 downto 0);
	signal addsub_carryout: std_logic;
	signal shift_result: std_logic_vector(31 downto 0);
	signal and_result: std_logic_vector(31 downto 0);
	signal or_result: std_logic_vector(31 downto 0);
	signal final_result: std_logic_vector(31 downto 0);

	-- ALU components	
	component adder_subtracter
		port(	datain_a: in std_logic_vector(31 downto 0);
			datain_b: in std_logic_vector(31 downto 0);
			add_sub: in std_logic;
			dataout: out std_logic_vector(31 downto 0);
			co: out std_logic);
	end component adder_subtracter;

	component shift_register
		port(	datain: in std_logic_vector(31 downto 0);
		   	dir: in std_logic;
			shamt:	in std_logic_vector(4 downto 0);
			dataout: out std_logic_vector(31 downto 0));
	end component shift_register;

begin
	-- Add ALU VHDL implementation here
	addsub: adder_subtracter port map(DataIn1, DataIn2, ALUCtrl(2), addsub_result, addsub_carryout);
	shift: shift_register port map(DataIn1, ALUCtrl(3), DataIn2(4 downto 0), shift_result);
	
	and_result <= DataIn1 and DataIn2;
	or_result <= DataIn1 or DataIn2;
	
	with ALUCtrl( 1 downto 0) select
		final_result <= addsub_result when "00",
				shift_result when "01",
				and_result when "10",
				or_result when others;

	with final_result select
		Zero <= '1' when  "00000000000000000000000000000000",
			'0' when others;

	ALUResult <= final_result;

end architecture ALU_Arch;



